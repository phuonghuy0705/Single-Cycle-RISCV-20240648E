module Instruction_Memory(rst,A,RD);

  input rst;
  input [31:0]A;
  output [31:0]RD;

  reg [31:0] mem [1023:0];
  
  assign RD = (~rst) ? {32{1'b0}} : mem[A[31:2]];

//   initial begin
//     $readmemh("memfile.hex",mem);
//   end



  initial begin  
    mem[0] = 32'h00028293;   //ADDI   0000_0000_0000_0010_1000_0010_1001_0011   //F3 -000 ->ADDI  // ADDI X5,X5,0  // X5 = 5 
    mem[1] = 32'h0062E233;   //OR     0000_0000_0110_0010_1110_0010_0011_0011   //F3 -110 ->OR    // OR X4,X5,X6   // X4 = 5 OR 4 = 5
    mem[2] = 32'h006273B3;   //AND    0000_0000_0110_0010_0111_0011_1011_0011   //F3 -111 ->AND   // AND X7,X4,X6  // X7 = 5 AND 4 = 4
    mem[3] = 32'h00638433;   //ADD    0000_0000_0110_0011_1000_0100_0011_0011   //F3 -000 ->ADD   // ADD X8,X7,X6  // X8 = 4 + 4 = 8
    mem[4] = 32'h404404B3;   //SUB    0100_0000_0100_0100_0000_0100_1011_0011   //F3 -000 ->SUB   // SUB X9,X8,X4  // X9 = 8 - 5 = 3
    mem[5] = 32'h0054C533;   //XOR    0000_0000_0101_0100_1100_0101_0011_0011   //F3 -100 ->XOR   // XOR X10,X9,X5 // X10 = 3 XOR 5 = 6
    mem[6] = 32'h0074A5B3;   //SLT    0000_0000_0111_0100_1010_0101_1011_0011   //F3 -010 ->SLT   // SLT X11,X9,X7 // X11 = 3 SLT 4 = 1
    mem[7] = 32'h0045A483;   //LW     0000_0000_0100_0101_1010_0100_1000_0011   //F3 -010 ->LW    // LW X9, 4(X11) // X9 = Mem[X11+4] = Mem[4]
    mem[8] = 32'h00752123;   //SW     0000_0000_0111_0101_0010_0001_0010_0011   //F3 -010 ->SW    // SW X7, 2(X10)  // Mem[X10+2] = Mem[8] = X7



  end

endmodule
