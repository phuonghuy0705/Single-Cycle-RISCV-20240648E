`timescale 1ns/1ps

module Register_File_tb;

    // Inputs
    reg clk, rst, WE3;
    reg [4:0] A1, A2, A3;
    reg [31:0] WD3;

    // Outputs
    wire [31:0] RD1, RD2;

    Register_File uut (
        .clk(clk),
        .rst(rst),
        .WE3(WE3),
        .WD3(WD3),
        .A1(A1),
        .A2(A2),
        .A3(A3),
        .RD1(RD1),
        .RD2(RD2)
    );

    always #5 clk = ~clk;

    initial begin

        clk = 0;
        rst = 0; WE3 = 0;
        A1 = 0; A2 = 0; A3 = 0; WD3 = 0;

        $display("==== Begin Register File Test ====");
        
        // Reset
        #10 rst = 1; // Turn on reset

        // Wait and check preloaded values
        #10;
        A1 = 5; A2 = 6;
        #10;
        $display("Read RD1 = R[5] = %d", RD1); // expect 5
        $display("Read RD2 = R[6] = %d", RD2); // expect 4

        // Test write to R[10]
        A3 = 10; WD3 = 32'h12345678; WE3 = 1;
        #10 WE3 = 0;

        // Read back from R[10]
        A1 = 10; A2 = 0;
        #10;
        $display("After write, R[10] = %h", RD1); // expect 0x12345678

        // Test write to R[0] (should not change)
        A3 = 0; WD3 = 32'hDEADBEEF; WE3 = 1;
        #10 WE3 = 0;

        A1 = 0;
        #10;
        $display("Attempted write to R[0], result = %h (should be 0)", RD1);

        $display("==== End of Test ====");
        $stop;
    end

endmodule

